-- $Id: $
-- File name:   rx_sr.vhd
-- Created:     9/29/2012
-- Author:      Vineeth Harikumar
-- Lab Section: 337-01
-- Version:     1.0  Initial Design Entry
-- Description: receiver shift register


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

entity rx_sr is
  port(
    clk : in std_logic;
    rst_n : in std_logic;
    sda_in : in std_logic;
    rising_edge_found : in std_logic;
    rx_enable : in std_logic;
    rx_data : out std_logic_vector(7 downto 0)
  );
end entity rx_sr;

architecture archRxSr of rx_sr is
	signal present_val : std_logic_vector(7 downto 0);
	signal next_val : std_logic_vector(7 downto 0);
  
begin
  
  REG: process (clk, rst_n)
  begin  -- process
		if('0' = rst_n) then
			present_val <= (others=>'0');
		elsif(rising_edge(clk)) then
			present_val <= next_val;
		end if; 
	end process;

	-- Next value logic: Shift in to the right when told to
	--next_val	<= sda_in & present_val(7 downto 1) when (('1' = rising_edge_found) and (rx_enable = '1') and rising_edge(clk)) else present_val;
	
	-- Output Logic
  rx_data	<= present_val(7 downto 0);
  
  nextValOutput : process(present_val, rising_edge_found, rx_enable)
  begin
    next_val <= present_val;
    if((rising_edge_found = '1') and (rx_enable = '1')) then
      --next_val <= sda_in & present_val(7 downto 1);
      next_val <= present_val(6 downto 0) & sda_in;
    end if;
  end process nextValOutput;
end architecture archRxSr;

